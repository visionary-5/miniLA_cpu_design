`timescale 1ns / 1ps
`include "defines.vh"

// ====================================================
// SEXT1 —— 立即数符号扩展单元1
// 支持 12位、16位、28位三种符号扩展类型
// 用于解析指令不同格式下的立即数
// ====================================================

// ===================================================
// ZEXT —— 零扩展单元
// 用于指令部分字段的无符号零扩展
// 常用于立即数的无符号型操作
// ===================================================

module EXIT_UNIT (
    input   wire [2:0]   sext1_op,     // 扩展类型选择
    input   wire [31:0]  inst,          // 原始指令

    output  wire [31:0]  sext1_ext,      // 扩展结果输出
    output  wire [31:0]  zext_ext       // 零扩展结果输出
);

    assign sext1_ext =
            (sext1_op == `EXT_OP_IMM12) ? {{20{inst[21]}}, inst[21:10]} :
            (sext1_op == `EXT_OP_IMM16) ? {{14{inst[25]}}, inst[25:10], 2'b0} :
            (sext1_op == `EXT_OP_IMM28) ? {{4{inst[9]}}, inst[9:0], inst[25:10], 2'b0} :
            32'b0;

    // 取指令第21~10位，前20位补零
    assign zext_ext = {20'b0, inst[21:10]};

endmodule   